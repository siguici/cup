module main

fn main() {
	println('👀 HTML/CSS inspired template rendering engine')
}
